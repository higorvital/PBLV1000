module Concertar_nome_3(
    input [11:0] wraddress_export,
    output [11:0] wraddress
);

    assign wraddress = wraddress_export;

endmodule