module Concertar_nome_2(
    input [11:0] rdaddress_export,
    output [11:0] rdaddress
);

    assign rdaddress = rdaddress_export;

endmodule